module Mux16(a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2, a1, a0, s, b);
   parameter k = 16;
   input [k-1:0] a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2, a1, a0;
   input [15:0]   s;
   output [k-1:0] b;
   assign b = (s[0]? a0 : 
        (s[1]? a1 :
         (s[2]? a2 :
          (s[3]? a3 :
           (s[4]? a4 :
            (s[5]? a5 :
             (s[6]? a6 :
			  (s[7]? a7 :
			   (s[8]? a8 :
			    (s[9]? a9 :
			     (s[10]? a10 :
			      (s[11]? a11 :
			       (s[12]? a12 :
			        (s[13]? a13 :
			         (s[14]? a14 : a15)))))))))))))));
endmodule // Mux16

module Mux32(a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2, a1, a0, s, b);
   parameter k = 32;
   input [k-1:0] a31, a30, a29, a28, a27, a26, a25, a24, a23, a22, a21, a20, 
					a19, a18, a17, a16, a15, a14, a13, a12, a11, a10, a9, a8, 
					a7, a6, a5, a4, a3, a2, a1, a0;
   input [15:0]   s;
   output [k-1:0] b;
   assign b = (s[0]? a0 : 
        (s[1]? a1 :
         (s[2]? a2 :
          (s[3]? a3 :
           (s[4]? a4 :
            (s[5]? a5 :
             (s[6]? a6 :
			  (s[7]? a7 :
			   (s[8]? a8 :
			    (s[9]? a9 :
			     (s[10]? a10 :
			      (s[11]? a11 :
			       (s[12]? a12 :
			        (s[13]? a13 :
			         (s[14]? a14 : a15)))))))))))))));
endmodule // Mux32

module testbench();
	reg [15:0] sel_16;
	reg [15:0] sel_32;
	reg [31:0] b15, b14, b13, b12, b11, b10, b9, b8, b7, b6, b5, b4, b3, b2, b1, b0;
	reg [15:0] a15;
	reg [15:0] a14;
	reg [15:0] a13;
	reg [15:0] a12;
	reg [15:0] a11;
	reg [15:0] a10;
	reg [15:0] a9;
	reg [15:0] a8;
	reg [15:0] a7;
	reg [15:0] a6;
	reg [15:0] a5;
	reg [15:0] a4;
	reg [15:0] a3;
	reg [15:0] a2;
	reg [15:0] a1;
	reg [15:0] a0;
	wire [15:0] aout;
	wire [31:0] bout;
	Mux16 mux0(a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2, 
					a1, a0, sel_16, aout);

	Mux32 mux1(b15, b14, b13, b12, b11, b10, b9, b8, b7, b6, 
							b5, b4, b3, b2, b1, b0, sel_32, bout);
	initial
		begin
		#10;
		sel_16 = 16'b0000000000000001;
		sel_32 = 16'b0000000000000010;
		a15 = 16'b1010101110101011;
      		a14 = 16'b0101011101010111;
                a13 = 16'b1010101110101011;
                a12 = 16'b0101011101010111;
		a11 = 16'b1010101110101011;
      		a10 = 16'b0101011101010111;
                a9 = 16'b1010101110101011;
                a8 = 16'b0101011101010111;
                a7 = 16'b1010101110101011;
                a6 = 16'b0101011101010111;
                a5 = 16'b1010101110101011;
                a4 = 16'b0101011101010111;
		a3 = 16'b0101011101010111;
                a2 = 16'b1010101110101011;
                a1 = 16'b0101011101010111;
                a0 = 16'b0101011101010000;
		b15 = 32'b10101011101010111010101110101011;
      		b14 = 32'b01010111010101110101011101010111;
                b13 = 32'b01010111010101110101011101010111;
                b12 = 32'b01010111010101110101011101010111;
		b11 = 32'b01010111010101110101011101010111;
      		b10 = 32'b01010111010101110101011101010111;
                b9 = 32'b01010111010101110101011101010111;
                b8 = 32'b01010111010101110101011101010111;
                b7 = 32'b01010111010101110101011101010111;
                b6 = 32'b01010111010101110101011101010111;
                b5 = 32'b01010111010101110101011101010111;
                b4 = 32'b01010111010101110101011101010111;
		b3 = 32'b01010111010101110101011101010111;
                b2 = 32'b01010111010101110101011101010111;
                b1 = 32'b01010111010101110101011101010000;
                b0 = 32'b01010111010101110101011101010111;
		$display(" Select for 32 bit is %b", sel_32);
		$display(" Select for 16 bit is %b", sel_16);
		#10;
		$display(" Value of of 32 bit 1st value is %b", b1);
		$display(" Value of of 16 bit 0th value is %b", a0);
		$display(" Value of mux32 is %b", bout);
		$display(" Value of mux16 is %b", aout);
	end
endmodule
