
module testbench();
initial begin
end
endmodule // testbench
